module clock_choice(

    input                       select,

    input                        latch,
    output                       s_clk,

	//////////// KEY //////////
	input 		     [1:0]		KEY
);

    


